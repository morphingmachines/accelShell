
module SimAccelTop #(
    // Width of hostCtrl data bus in bits
    parameter HOSTCTRL_DATA_WIDTH = 32,
    // Width of hostCtrl address bus in bits
    parameter HOSTCTRL_ADDR_WIDTH = 16,
    // Width of hostCtrl wstrb 
    parameter HOSTCTRL_STRB_WIDTH = (HOSTCTRL_DATA_WIDTH / 8),
    // Width of hostCtrl ID signal
    parameter HOSTCTRL_ID_WIDTH = 8,
    // Width of dma data bus in bits
    parameter HOSTMEM_DATA_WIDTH = 32,
    // Width of dma address bus in bits
    parameter HOSTMEM_ADDR_WIDTH = 16,
    // Width of dma wstrb 
    parameter HOSTMEM_STRB_WIDTH = (HOSTMEM_DATA_WIDTH / 8),
    // Width of dma ID signal
    parameter HOSTMEM_ID_WIDTH = 8
) (
    input wire clk,
    input wire rst,

    output wire                           hostCtrl_awready,
    input  wire                           hostCtrl_awvalid,
    input  wire [  HOSTCTRL_ID_WIDTH-1:0] hostCtrl_awid,
    input  wire [HOSTCTRL_ADDR_WIDTH-1:0] hostCtrl_awaddr,
    input  wire [                    7:0] hostCtrl_awlen,
    input  wire [                    2:0] hostCtrl_awsize,
    input  wire [                    1:0] hostCtrl_awburst,
    input  wire                           hostCtrl_awlock,
    input  wire [                    3:0] hostCtrl_awcache,
    input  wire [                    2:0] hostCtrl_awprot,
    output wire                           hostCtrl_wready,
    input  wire                           hostCtrl_wvalid,
    input  wire [HOSTCTRL_DATA_WIDTH-1:0] hostCtrl_wdata,
    input  wire [HOSTCTRL_STRB_WIDTH-1:0] hostCtrl_wstrb,
    input  wire                           hostCtrl_wlast,
    input  wire                           hostCtrl_bready,
    output wire                           hostCtrl_bvalid,
    output wire [  HOSTCTRL_ID_WIDTH-1:0] hostCtrl_bid,
    output wire [                    1:0] hostCtrl_bresp,
    output wire                           hostCtrl_arready,
    input  wire                           hostCtrl_arvalid,
    input  wire [  HOSTCTRL_ID_WIDTH-1:0] hostCtrl_arid,
    input  wire [HOSTCTRL_ADDR_WIDTH-1:0] hostCtrl_araddr,
    input  wire [                    7:0] hostCtrl_arlen,
    input  wire [                    2:0] hostCtrl_arsize,
    input  wire [                    1:0] hostCtrl_arburst,
    input  wire                           hostCtrl_arlock,
    input  wire [                    3:0] hostCtrl_arcache,
    input  wire [                    2:0] hostCtrl_arprot,
    input  wire                           hostCtrl_rready,
    output wire                           hostCtrl_rvalid,
    output wire [  HOSTCTRL_ID_WIDTH-1:0] hostCtrl_rid,
    output wire [HOSTCTRL_DATA_WIDTH-1:0] hostCtrl_rdata,
    output wire [                    1:0] hostCtrl_rresp,
    output wire                           hostCtrl_rlast,
    output wire                           hostMem_awready,
    input  wire                           hostMem_awvalid,
    input  wire [   HOSTMEM_ID_WIDTH-1:0] hostMem_awid,
    input  wire [ HOSTMEM_ADDR_WIDTH-1:0] hostMem_awaddr,
    input  wire [                    7:0] hostMem_awlen,
    input  wire [                    2:0] hostMem_awsize,
    input  wire [                    1:0] hostMem_awburst,
    input  wire                           hostMem_awlock,
    input  wire [                    3:0] hostMem_awcache,
    input  wire [                    2:0] hostMem_awprot,
    output wire                           hostMem_wready,
    input  wire                           hostMem_wvalid,
    input  wire [ HOSTMEM_DATA_WIDTH-1:0] hostMem_wdata,
    input  wire [ HOSTMEM_STRB_WIDTH-1:0] hostMem_wstrb,
    input  wire                           hostMem_wlast,
    input  wire                           hostMem_bready,
    output wire                           hostMem_bvalid,
    output wire [   HOSTMEM_ID_WIDTH-1:0] hostMem_bid,
    output wire [                    1:0] hostMem_bresp,
    output wire                           hostMem_arready,
    input  wire                           hostMem_arvalid,
    input  wire [   HOSTMEM_ID_WIDTH-1:0] hostMem_arid,
    input  wire [ HOSTMEM_ADDR_WIDTH-1:0] hostMem_araddr,
    input  wire [                    7:0] hostMem_arlen,
    input  wire [                    2:0] hostMem_arsize,
    input  wire [                    1:0] hostMem_arburst,
    input  wire                           hostMem_arlock,
    input  wire [                    3:0] hostMem_arcache,
    input  wire [                    2:0] hostMem_arprot,
    input  wire                           hostMem_rready,
    output wire                           hostMem_rvalid,
    output wire [   HOSTMEM_ID_WIDTH-1:0] hostMem_rid,
    output wire [ HOSTMEM_DATA_WIDTH-1:0] hostMem_rdata,
    output wire [                    1:0] hostMem_rresp,
    output wire                           hostMem_rlast
);

  SimAccel simAccel (
      .clock(clk),
      .reset(rst),
      .hostCtrl_0_aw_ready(hostCtrl_awready),
      .hostCtrl_0_aw_valid(hostCtrl_awvalid),
      .hostCtrl_0_aw_bits_id(hostCtrl_awid),
      .hostCtrl_0_aw_bits_addr(hostCtrl_awaddr),
      .hostCtrl_0_aw_bits_len(hostCtrl_awlen),
      .hostCtrl_0_aw_bits_size(hostCtrl_awsize),
      .hostCtrl_0_aw_bits_burst(hostCtrl_awburst),
      .hostCtrl_0_aw_bits_lock(hostCtrl_awlock),
      .hostCtrl_0_aw_bits_cache(hostCtrl_awcache),
      .hostCtrl_0_aw_bits_prot(hostCtrl_awprot),
      .hostCtrl_0_aw_bits_qos(3'b0),
      .hostCtrl_0_w_ready(hostCtrl_wready),
      .hostCtrl_0_w_valid(hostCtrl_wvalid),
      .hostCtrl_0_w_bits_data(hostCtrl_wdata),
      .hostCtrl_0_w_bits_strb(hostCtrl_wstrb),
      .hostCtrl_0_w_bits_last(hostCtrl_wlast),
      .hostCtrl_0_b_ready(hostCtrl_bready),
      .hostCtrl_0_b_valid(hostCtrl_bvalid),
      .hostCtrl_0_b_bits_id(hostCtrl_bid),
      .hostCtrl_0_b_bits_resp(hostCtrl_bresp),
      .hostCtrl_0_ar_ready(hostCtrl_arready),
      .hostCtrl_0_ar_valid(hostCtrl_arvalid),
      .hostCtrl_0_ar_bits_id(hostCtrl_arid),
      .hostCtrl_0_ar_bits_addr(hostCtrl_araddr),
      .hostCtrl_0_ar_bits_len(hostCtrl_arlen),
      .hostCtrl_0_ar_bits_size(hostCtrl_arsize),
      .hostCtrl_0_ar_bits_burst(hostCtrl_arburst),
      .hostCtrl_0_ar_bits_lock(hostCtrl_arlock),
      .hostCtrl_0_ar_bits_cache(hostCtrl_arcache),
      .hostCtrl_0_ar_bits_prot(hostCtrl_arprot),
      .hostCtrl_0_ar_bits_qos(3'b0),
      .hostCtrl_0_r_ready(hostCtrl_rready),
      .hostCtrl_0_r_valid(hostCtrl_rvalid),
      .hostCtrl_0_r_bits_id(hostCtrl_rid),
      .hostCtrl_0_r_bits_data(hostCtrl_rdata),
      .hostCtrl_0_r_bits_resp(hostCtrl_rresp),
      .hostCtrl_0_r_bits_last(hostCtrl_rlast),
      .hostMem_0_aw_ready(hostMem_awready),
      .hostMem_0_aw_valid(hostMem_awvalid),
      .hostMem_0_aw_bits_id(hostMem_awid),
      .hostMem_0_aw_bits_addr(hostMem_awaddr),
      .hostMem_0_aw_bits_len(hostMem_awlen),
      .hostMem_0_aw_bits_size(hostMem_awsize),
      .hostMem_0_aw_bits_burst(hostMem_awburst),
      .hostMem_0_aw_bits_lock(hostMem_awlock),
      .hostMem_0_aw_bits_cache(hostMem_awcache),
      .hostMem_0_aw_bits_prot(hostMem_awprot),
      .hostMem_0_aw_bits_qos(3'b0),
      .hostMem_0_w_ready(hostMem_wready),
      .hostMem_0_w_valid(hostMem_wvalid),
      .hostMem_0_w_bits_data(hostMem_wdata),
      .hostMem_0_w_bits_strb(hostMem_wstrb),
      .hostMem_0_w_bits_last(hostMem_wlast),
      .hostMem_0_b_ready(hostMem_bready),
      .hostMem_0_b_valid(hostMem_bvalid),
      .hostMem_0_b_bits_id(hostMem_bid),
      .hostMem_0_b_bits_resp(hostMem_bresp),
      .hostMem_0_ar_ready(hostMem_arready),
      .hostMem_0_ar_valid(hostMem_arvalid),
      .hostMem_0_ar_bits_id(hostMem_arid),
      .hostMem_0_ar_bits_addr(hostMem_araddr),
      .hostMem_0_ar_bits_len(hostMem_arlen),
      .hostMem_0_ar_bits_size(hostMem_arsize),
      .hostMem_0_ar_bits_burst(hostMem_arburst),
      .hostMem_0_ar_bits_lock(hostMem_arlock),
      .hostMem_0_ar_bits_cache(hostMem_arcache),
      .hostMem_0_ar_bits_prot(hostMem_arprot),
      .hostMem_0_ar_bits_qos(3'b0),
      .hostMem_0_r_ready(hostMem_rready),
      .hostMem_0_r_valid(hostMem_rvalid),
      .hostMem_0_r_bits_id(hostMem_rid),
      .hostMem_0_r_bits_data(hostMem_rdata),
      .hostMem_0_r_bits_resp(hostMem_rresp),
      .hostMem_0_r_bits_last(hostMem_rlast),
      .io_accelDomain_clock(clk),
      .io_accelDomain_reset(rst)
  );
endmodule
