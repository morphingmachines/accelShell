
module SimDeviceMemTop #(
    // Width of dma data bus in bits
    parameter HOSTMEM_DATA_WIDTH = 32,
    // Width of dma address bus in bits
    parameter HOSTMEM_ADDR_WIDTH = 16,
    // Width of dma wstrb 
    parameter HOSTMEM_STRB_WIDTH = (HOSTMEM_DATA_WIDTH / 8),
    // Width of dma ID signal
    parameter HOSTMEM_ID_WIDTH   = 8
) (
    input wire clk,
    input wire rst,

    output wire                          hostMem_awready,
    input  wire                          hostMem_awvalid,
    input  wire [  HOSTMEM_ID_WIDTH-1:0] hostMem_awid,
    input  wire [HOSTMEM_ADDR_WIDTH-1:0] hostMem_awaddr,
    input  wire [                   7:0] hostMem_awlen,
    input  wire [                   2:0] hostMem_awsize,
    input  wire [                   1:0] hostMem_awburst,
    input  wire                          hostMem_awlock,
    input  wire [                   3:0] hostMem_awcache,
    input  wire [                   2:0] hostMem_awprot,
    output wire                          hostMem_wready,
    input  wire                          hostMem_wvalid,
    input  wire [HOSTMEM_DATA_WIDTH-1:0] hostMem_wdata,
    input  wire [HOSTMEM_STRB_WIDTH-1:0] hostMem_wstrb,
    input  wire                          hostMem_wlast,
    input  wire                          hostMem_bready,
    output wire                          hostMem_bvalid,
    output wire [  HOSTMEM_ID_WIDTH-1:0] hostMem_bid,
    output wire [                   1:0] hostMem_bresp,
    output wire                          hostMem_arready,
    input  wire                          hostMem_arvalid,
    input  wire [  HOSTMEM_ID_WIDTH-1:0] hostMem_arid,
    input  wire [HOSTMEM_ADDR_WIDTH-1:0] hostMem_araddr,
    input  wire [                   7:0] hostMem_arlen,
    input  wire [                   2:0] hostMem_arsize,
    input  wire [                   1:0] hostMem_arburst,
    input  wire                          hostMem_arlock,
    input  wire [                   3:0] hostMem_arcache,
    input  wire [                   2:0] hostMem_arprot,
    input  wire                          hostMem_rready,
    output wire                          hostMem_rvalid,
    output wire [  HOSTMEM_ID_WIDTH-1:0] hostMem_rid,
    output wire [HOSTMEM_DATA_WIDTH-1:0] hostMem_rdata,
    output wire [                   1:0] hostMem_rresp,
    output wire                          hostMem_rlast
);

  SimDeviceMem simDeviceMem (
      .clock(clk),
      .reset(rst),
      .hostMem_0_aw_ready(hostMem_awready),
      .hostMem_0_aw_valid(hostMem_awvalid),
      .hostMem_0_aw_bits_id(hostMem_awid),
      .hostMem_0_aw_bits_addr(hostMem_awaddr),
      .hostMem_0_aw_bits_len(hostMem_awlen),
      .hostMem_0_aw_bits_size(hostMem_awsize),
      .hostMem_0_aw_bits_burst(hostMem_awburst),
      .hostMem_0_aw_bits_lock(hostMem_awlock),
      .hostMem_0_aw_bits_cache(hostMem_awcache),
      .hostMem_0_aw_bits_prot(hostMem_awprot),
      .hostMem_0_aw_bits_qos(3'b0),
      .hostMem_0_w_ready(hostMem_wready),
      .hostMem_0_w_valid(hostMem_wvalid),
      .hostMem_0_w_bits_data(hostMem_wdata),
      .hostMem_0_w_bits_strb(hostMem_wstrb),
      .hostMem_0_w_bits_last(hostMem_wlast),
      .hostMem_0_b_ready(hostMem_bready),
      .hostMem_0_b_valid(hostMem_bvalid),
      .hostMem_0_b_bits_id(hostMem_bid),
      .hostMem_0_b_bits_resp(hostMem_bresp),
      .hostMem_0_ar_ready(hostMem_arready),
      .hostMem_0_ar_valid(hostMem_arvalid),
      .hostMem_0_ar_bits_id(hostMem_arid),
      .hostMem_0_ar_bits_addr(hostMem_araddr),
      .hostMem_0_ar_bits_len(hostMem_arlen),
      .hostMem_0_ar_bits_size(hostMem_arsize),
      .hostMem_0_ar_bits_burst(hostMem_arburst),
      .hostMem_0_ar_bits_lock(hostMem_arlock),
      .hostMem_0_ar_bits_cache(hostMem_arcache),
      .hostMem_0_ar_bits_prot(hostMem_arprot),
      .hostMem_0_ar_bits_qos(3'b0),
      .hostMem_0_r_ready(hostMem_rready),
      .hostMem_0_r_valid(hostMem_rvalid),
      .hostMem_0_r_bits_id(hostMem_rid),
      .hostMem_0_r_bits_data(hostMem_rdata),
      .hostMem_0_r_bits_resp(hostMem_rresp),
      .hostMem_0_r_bits_last(hostMem_rlast)
  );
endmodule
